-- test 

