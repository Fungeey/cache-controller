library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity CacheController is
	Port    (	clk 				: in  STD_LOGIC;
				reset				
				addr_in			: in 	STD_LOGIC_VECTOR(15 downto 0));
end CacheController;
